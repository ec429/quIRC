int:width:80:30:::width:width:S:display width
int:height:24:5:::height:height:S:display height
int:mirc_colour_compat:1:0:2:mcc:mcc:mcc:L:mirc colour compatibility
int:force_redraw:0:0:3:fred:fred:fred:L:force-redraw
int:buflines:1024:32::buf:buf-lines:buf:S:buffer lines
int:maxnlen:16:4::mnln:maxnicklen:mnln:S:max nick length
bool:full_width_colour:false:::fwc:fwc:fwc:B:full width colour
bool:hilite_tabstrip:false:::hts:hts:hts:B:highlight tabstrip
bool:tsb:true:::tsb:tsb:tsb:B:top status bar
int:tping:30:15::tping:tping:tping:S:outbound ping time
int:ts:1:0:4:ts:timestamps:ts:L:timestamping
bool:utc:false:::utc:utc:utc:B:UTC timestamps
bool:its:false:::its:its:its:B:input clock
bool:quiet:false:::quiet:quiet:quiet:B:quiet mode
bool:debug:false:::debug:debug:debug:B:debugging
bool:conf:false:::conf:conf::B:conference mode (default)
bool:show_prefix:false:::prefix:prefix:prefix:B:display nick prefixes
bool:titles:true:::titles:titles:titles:B:xterm title
bool:winch:true:::winch:winch:winch:B:react to SIGWINCH (window change)
